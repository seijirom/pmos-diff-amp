**.subckt currentsource_test14umWilson Vout Vout2 Vout
*.opin Vout
*.opin Vout2
*.opin Vout
V1 GND net8 5
M1 net3 net3 net1 net1 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=20
V2 net1 GND 5
I1 net6 net8 200u
M2 net5 net3 net1 net1 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=20
V3 Vout GND 5
M3 net6 net6 net5 net1 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=40
M4 Vout net6 net3 net1 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=40
V4 GND net9 5
M5 net4 net4 net2 net2 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=30
V5 net2 GND 5
I2 net7 net9 200u
M6 net7 net4 net2 net2 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=30
M8 Vout2 net7 net4 net2 YSS_PMOS w=14u l=14u as=0 ps=0 ad=0 pd=0 m=40
E1 Vout2 GND Vout GND 1.0
**** begin user architecture code

.include ../parameter2/mineda2020_1_pmos.txt


.dc V3 -5 5 20m

**** end user architecture code
**.ends
.GLOBAL GND
.end
